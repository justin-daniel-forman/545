`define NOP 8'h00
`define INC 8'b00???100
