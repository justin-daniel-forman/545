//-----------------------------------------------------------------------------
//datapath
//  This module contains the main datapath for the system. It operates on 
//  a shared internal databus that can drive the external data bus. Only 
//  one component from the datapath can drive the databus at a given time.
//-----------------------------------------------------------------------------
module datapath (


);

endmodule: datapath
