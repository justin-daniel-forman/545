module psg_top (

  //---------------------------------------------------------------------------
  //Bus Interface
  //  - data_bus:
  //  - addr_bus:
  //---------------------------------------------------------------------------
  inout wire [7:0]   data_bus,
  inout wire [15:0]  addr_bus,


  //---------------------------------------------------------------------------
  //Board output interface
  //
  //---------------------------------------------------------------------------

);



endmodule: psg_top
