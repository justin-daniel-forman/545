`define NOP 8'h00
`define INC 8'b00???100

`define EXT_INST 8'hED
`define LDI      8'hA0


//ALU commands
`define INCR_A  4'b0001
`define DECR_A  4'b0010
`define ALU_NOP 4'b0000
