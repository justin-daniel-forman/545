`define NOP 8'h00
`define INC 8'b00???100


//ALU commands
`define INCR_A 4'b0001
