`define NOP 8'h00
`define INC 8'b00???100

`define INC_IX_0 8'hDD
`define INC_IX_1 8'h23

//ALU commands
`define INCR_A  4'b0001
`define ALU_NOP 4'b0000
